// full adder using half adder 

module rpa(input a,b,cin ,output sum,cout);
 
  FA_using_HA add1(a,b,cin,sum,cout);

endmodule