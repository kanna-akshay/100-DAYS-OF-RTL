// ripple carry subractor 

module rps(input a,b,Bout ,output diff,Bin);
 
  FS_using_HS diff1(a,b,Bout,diff,Bin);

endmodule